library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_textio.all;  -- For logic types I/O
library std;
use IEEE.numeric_std.all;
use std.env.all;                -- For hierarchical/external signals
use std.textio.all;             -- For basic I/O


entity tb_proj2_hardware_regs is 
    generic (gClk_per: time:= 10ns; N : integer := 32);
end entity;

architecture tb_arch_proj2_hardware_regs of tb_proj2_hardware_regs is
--components

--signals

--begin

begin

end tb_arch_proj2_hardware_regs ; -- tb_arch_proj2_hardware_regs
